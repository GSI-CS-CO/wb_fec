library verilog;
use verilog.vl_types.all;
entity main is
end main;
