library verilog;
use verilog.vl_types.all;
entity main_sv_unit is
end main_sv_unit;
